`ifndef APB_TESTS_SVH
`define APB_TESTS_SVH

`include "apb_base_test.sv"

// apb3 tests
`include "apb3_single_trans_test.sv"
`include "apb3_burst_trans_test.sv"

// apb4 tests
`include "apb4_single_trans_test.sv"

`endif