`ifndef APB_SEQUENCES_SVH
`define APB_SEQUENCES_SVH

`include "apb_base_virtual_sequence.sv"

// apb3 virt seq
`include "apb3_single_trans_virt_seq.sv"
`include "apb3_burst_trans_virt_seq.sv"

// apb4 virt seq
`include "apb4_single_trans_virt_seq.sv"

`endif